module inversora //definindo o módulo
(
	input in,
	output out
);

assign out = ~in;
endmodule
 